package pb_pkg;

  `include "inter.sv"
  `include "trans.sv"
  `include "gens.sv"
  `include "dr.sv"
  `include "mo.sv"
  `include "sc.sv"
  `include "en.sv"
  `include "tes.sv"

endpackage
